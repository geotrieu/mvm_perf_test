// static_params.vh

`ifndef _static_params_vh_
`define _static_params_vh_

`define DATAW 64
`define FIFO_DEPTH 8

`define AXIS_IDW 2
`define AXIS_DESTW 4
`define AXIS_MAX_DATAW 64

`endif //_static_params_vh_
