// config.vh

`ifndef _config_vh_
`define _config_vh_

`define PROJECT_DIR "/home/gtrieu/projects/mvm_perf_test/noc/"

`endif //_config_vh_
