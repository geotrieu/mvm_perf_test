// config.vh

`ifndef _config_vh_
`define _config_vh_

`define PROJECT_DIR "~/projects/mvm_perf_test/noc/sim"

`endif //_config_vh_
